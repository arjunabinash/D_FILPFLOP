interface dff_if;
  logic din;
  logic dout;
  logic rst;
  logic clk;
endinterface